module mod_a (
    input in1, in2,
    output out
    );

endmodule
