// A Module can contain instances of other modules 
// And this is how a larger complex circuits are designed 

module mod_a (
    input in1, in2,
    output out,
    );

endmodule


module top_module (
    input a,b,
    output out
    );

    
endmodule